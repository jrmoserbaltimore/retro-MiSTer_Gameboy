// vim: sw=4 ts=4 et
// Copyright (c) 2020 Moonset Technologies, LLC
// License:  MIT, see LICENSE.md
//
// Game Boy Color Shim.  The shim sets up for an actual core, creating RAM objects, mapping the
// expansion port (e.g. to a cartridge), exposing the controller properly to the core, managing
// CATC, handling cache, and so forth.

// This is the core shim.  RetroConosle connects everything to this, which then connects to the
// core module.  In here we set up various types of RAM, clock control, the cartridge controller,
// and any peripherals.
//
// Detecting DMG, CGB, GBA:
//   - DMG:  CPU A register == 0x01 (also SGB)
//   - MGB:  CPU A register == 0xff (Gameboy Pocket, SGB2)
//   - CGB:  CPU A register == 0x11, B[0] == 0
//   - GBA:  CPU A register == 0x11, B[0] == 1 
module RetroCoreShim
#(
    parameter DeviceType = "Xilinx",
    parameter CoreClock = 200000000 // 200MHz FPGA core clock
)
(
    // The console sends a core system clock (e.g. 200MHz) to produce the reference clock.
    ISysCon SysCon, // Core system clock

    // DDR System RAM or other large RAM.

    IWishbone.Initiator MainRAM,
    // DDR, HyperRAM, or SRAM on the expansion bus
    IWishbone.Initiator ExpansionRAM0,
    IWishbone.Initiator ExpansionRAM1,
    IWishbone.Initiator ExpansionRAM2,

    output logic [23:0] Video,
    output logic [23:0] Audio, // 96kHz 24-bit, downsample to 48kHz 16-bit
    // ================
    // = External Bus =
    // ================

    // Cartridge bus wide enough for NES, 69 I/O
    output logic CartridgeClk,
//    input logic [68:0] CartridgeIn,
//    output logic [68:0] CartridgeOut,

    // Controller I/O, from �C
    input logic ControllerIn,
    output logic ControllerOut,

    // Expansion
    input logic [31:0] ExpansionPortIn,
    output logic [31:0] ExpansionPortOut,

    // Console
    IWishbone.Target Host
);

    wire Delay;
    wire Reset;
    wire Ce;
    
    wire Read, Write;
    wire [15:0] Address;
    wire [7:0] DataIn, DataOut;
    wire AudioIn;
    wire CS, Ready, DataReady;

    wire CartDelay;
    wire MainRAMDelay;
    wire VRAMDelay;
    
    // The cartridge controller needs to always provide both Ready and DataReady unless waiting
    // for operations.  These may frequently fall between clock ticks.  When using a hardware
    // cartridge, both of these should be kept on.
    assign Delay = ~(Ready & DataReady);

    // ======================
    // = System RAM Objects =
    // ======================
    // We create BRAMs in the shim so a different shim can use the GBC Cartridge Controller without
    // dedicating the BRAM exclusively to the GBC when not running.
    IWishbone
    #(
        .AddressWidth(15),
        .DataWidth(8) 
    ) IGBSystemRAM();

    //(* dont_touch = "true" *)
    WishboneBRAM
    #(
        .AddressWidth(15),
        .DataWidth(8),
        .DeviceType(DeviceType)
    ) GBSystemRAM
    (
        .SysCon(SysCon),
        .Initiator(IGBSystemRAM.Target)
    );

    IWishbone
    #(
        .AddressWidth(14),
        .DataWidth(8) 
    ) IGBVideoRAM();

    //(* dont_touch = "true" *)
    WishboneBRAM
    #(
        .AddressWidth(14),
        .DataWidth(8),
        .DeviceType(DeviceType)
    ) GBVideoRAM
    (
        .SysCon(SysCon),
        .Initiator(IGBVideoRAM.Target)
    );
    
    IWishbone
    #(
        .AddressWidth(17),
        .DataWidth(8) 
    ) IGBCartridgeRAM();

    //(* dont_touch = "true" *)
    WishboneBRAM
    #(
        .AddressWidth(17),
        .DataWidth(8),
        .DeviceType(DeviceType)
    ) GBCartridgeRAM
    (
        .SysCon(SysCon),
        .Initiator(IGBCartridgeRAM.Target)
    );
    // TODO:  Chunk of BRAM for cartridge cache
    // TODO:  Chunk of BRAM for mappers

    // ========
    // = CATC =
    // ========
    // Cartridge controller triggers Delay if data isn't ready
    /*
    RetroCATC CATC(
        .Clk(CoreClk),
        .Delay(Delay),
        .ClkEn(ClkEn),
        .Reset(Reset),
        .ClkEnOut(Ce)
    );
    */

    // =================================
    // = Interface to hardware GamePak =
    // =================================
    /*
    IGBCGamePak GamePak(
        .Clk(CartridgeClk),
        .Write(CartridgeOut[2]),
        .Read(CartridgeOut[3]),
        .CS(CartridgeOut[4]),
        .Address(CartridgeOut[20:5]),
        .DFromPak(CartridgeIn[28:21]),
        .DToPak(CartridgeOut[28:21]),
        .Reset(CartridgeOut[29]),
        .Audio(CartridgeIn[30])
    );
    */

    // ========================
    // = Interface to GamePak =
    // ========================

    IWishbone
    #(
        .AddressWidth(16),
        .DataWidth(8)
    )
    ISystemBus();

    IWishbone
    #(
        .AddressWidth(16),
        .DataWidth(8)
    )
    IRTC();
    // FIXME:  Hastily-assembled stuff to get this to actually synthesize
    
    IWishbone
    #(
        .AddressWidth(23),
        .DataWidth(8) 
    ) ILoadImage();

    // XXX:  Need to instantiate a cache here, not an 8MB BRAM
    //(* dont_touch = "true" *)
    /*
    WishboneBRAM
    #(
        .AddressWidth(23),
        .DataWidth(8),
        .DeviceType(DeviceType)
    ) LoadImage
    (
        .SysCon(SysCon),
        .Initiator(ILoadImage.Target)
    );
    */
    IWishbone
    #(
        .AddressWidth(16),
        .DataWidth(8)
    )
    IMapper();

    //(* dont_touch = "true" *)
    GBCMapper Mapper
    (
        .SysCon(SysCon),
        //.LoadImage(ILoadImage.Initiator),
        .LoadImage(ExpansionRAM0),
        .CartridgeRAM(IGBCartridgeRAM.Initiator),
        .RTC(IRTC.Initiator), // XXX:  Placeholder
        .MemoryBus(IMapper.Target)
    );

    //(* dont_touch = "true" *)
    GBCMemoryBus SystemBus
    (
        .SysCon(SysCon),
        // System and video BRAMs
        .SystemRAM(IGBSystemRAM.Initiator),
        .VideoRAM(IGBVideoRAM.Initiator),
        .VideoStatus(3'b000),
        .Cartridge(IMapper.Initiator),
        .MemoryBus(Host) // Placeholder 
    );

    logic [15:0] addrct;
    
    always_ff @(posedge SysCon.CLK)
    begin
        if (SysCon.RST)
        begin
            Host.Unstall();
        end
    end
    /*
    RetroMyCore TheCore
    (
        .Clk(CoreClk),
        .ClkEn(Ce),
        .AV(AV),
        .MemoryBus(GamePakFrontend.Initiator),
        .GamePak(GamePakBus.Gameboy),
        // TODO:  Serial controller
        // etc.
        .SerialOut(0),
        .SerialIn(0),
        .SD(0),
        .SerialClk(0)
    );
    */
endmodule